
module spi_node (
    
);
    
endmodule